// Opcode
`define OPCODE_R        7'b0110011
`define OPCODE_I        7'b0010011
`define OPCODE_LW       7'b0000011
`define OPCODE_JALR     7'b1100111
`define OPCODE_SW       7'b0100011
`define OPCODE_B        7'b1100011
`define OPCODE_LUI      7'b0110111
`define OPCODE_JAL      7'b1101111
